`timescale 1ns / 1ps
//Author: Murat Celik
//Date : 02.09.2023
//N=16 Mux
//Test Bench


module n1_mux_tb;
	reg [15:0] in;
	reg [3:0] sel;
	wire y;
	//UUT
	n1_mux uut (
		.in(in), 
		.sel(sel), 
		.y(y)
	);
//Tests
initial begin
in=16'b1000000000000000; sel=4'b0000; 
#10 in=16'b0100000000000010; sel=4'b0001; 
#10 in=16'b0010000000000100; sel=4'b0010;
#10 in=16'b0001000000000000; sel=4'b0011;
#10 in=16'b0000100000011000; sel=4'b0100; 
#10 in=16'b0000010000000000; sel=4'b0101; 
#10 in=16'b0000001000000000; sel=4'b0110;
#10 in=16'b0000000111100000; sel=4'b0111;
#10 in=16'b0000000010000000; sel=4'b1000;
#10 in=16'b0000000001000000; sel=4'b1001;
#10 in=16'b0000011000100000; sel=4'b1010; 
#10 in=16'b0000000000010000; sel=4'b1011;
#10 in=16'b0000000000001000; sel=4'b1100; 
#10 in=16'b0000000000000100; sel=4'b1101; 
#10 in=16'b0000000000000010; sel=4'b1110; 
#10 in=16'b1000000000000001; sel=4'b1111;
end 
initial
begin
$monitor("in=%b | sel=%b | out=%b",in,sel,y);			 
#500 $finish;
end     
endmodule
